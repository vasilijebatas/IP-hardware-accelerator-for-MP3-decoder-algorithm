----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08/08/2023 11:19:02 AM
-- Design Name: 
-- Module Name: rom_lut - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with ununsigned or ununsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_cos is
Generic(
        WIDTH_D: positive;
        WIDTH_A: positive;
        DEPTH: positive
    );
    Port (
        clk: in std_logic;

        angle: in std_logic_vector(WIDTH_A-1 downto 0);
        cos: out std_logic_vector(WIDTH_D-1 downto 0);

        en: in std_logic
    );
end rom_cos;

architecture syn of rom_cos is
    
    
    
    type rom_type is array(0 to DEPTH-1) of std_logic_vector(WIDTH_D-1 downto 0);
    signal ROM: rom_type :=(
        "0100000000000000", 
        "0011111111111101", 
        "0011111111110110", 
        "0011111111101001", 
        "0011111111011000", 
        "0011111111000001", 
        "0011111110100110", 
        "0011111110000110", 
        "0011111101100000", 
        "0011111100110110", 
        "0011111100000111", 
        "0011111011010011", 
        "0011111010011010", 
        "0011111001011100", 
        "0011111000011001", 
        "0011110111010010", 
        "0011110110000101", 
        "0011110100110100", 
        "0011110011011110", 
        "0011110010000100", 
        "0011110000100100", 
        "0011101111000000", 
        "0011101101011000", 
        "0011101011101010", 
        "0011101001111000", 
        "0011101000000010", 
        "0011100110000111", 
        "0011100100001000", 
        "0011100010000100", 
        "0011011111111011", 
        "0011011101101111", 
        "0011011011011110", 
        "0011011001001000", 
        "0011010110101111", 
        "0011010100010001", 
        "0011010001101111", 
        "0011001111001010", 
        "0011001100100000", 
        "0011001001110010", 
        "0011000111000000", 
        "0011000100001010", 
        "0011000001010001", 
        "0010111110010011", 
        "0010111011010010", 
        "0010111000001110", 
        "0010110101000101", 
        "0010110001111010", 
        "0010101110101010", 
        "0010101011011000", 
        "0010101000000010", 
        "0010100100101000", 
        "0010100001001100", 
        "0010011101101100", 
        "0010011010001010", 
        "0010010110100100", 
        "0010010010111100", 
        "0010001111010000", 
        "0010001011100010", 
        "0010000111110001", 
        "0010000011111101", 
        "0010000000000111", 
        "0001111100001110", 
        "0001111000010011", 
        "0001110100010110", 
        "0001110000010110", 
        "0001101100010100", 
        "0001101000010000", 
        "0001100100001010", 
        "0001100000000010", 
        "0001011011111000", 
        "0001010111101101", 
        "0001010011011111", 
        "0001001111010000", 
        "0001001011000000", 
        "0001000110101110", 
        "0001000010011010", 
        "0000111110000110", 
        "0000111001110000", 
        "0000110101011001", 
        "0000110001000001", 
        "0000101100101000", 
        "0000101000001110", 
        "0000100011110011", 
        "0000011111011000", 
        "0000011010111100", 
        "0000010110100000", 
        "0000010010000011", 
        "0000001101100110", 
        "0000001001001000", 
        "0000000100101010", 
        "0000000000001101", 
        "0000000100010000", 
        "0000001000101110", 
        "0000001101001100", 
        "0000010001101001", 
        "0000010110000110", 
        "0000011010100010", 
        "0000011110111110", 
        "0000100011011010", 
        "0000100111110100", 
        "0000101100001110", 
        "0000110000100111", 
        "0000110100111111", 
        "0000111001010111", 
        "0000111101101101", 
        "0001000010000001", 
        "0001000110010101", 
        "0001001010100111", 
        "0001001110111000", 
        "0001010011000111", 
        "0001010111010100", 
        "0001011011100000", 
        "0001011111101010", 
        "0001100011110010", 
        "0001100111111000", 
        "0001101011111101", 
        "0001101111111111", 
        "0001110011111111", 
        "0001110111111100", 
        "0001111011111000", 
        "0001111111110000", 
        "0010000011100111", 
        "0010000111011011", 
        "0010001011001100", 
        "0010001110111010", 
        "0010010010100110", 
        "0010010110001111", 
        "0010011001110101", 
        "0010011101011000", 
        "0010100000111000", 
        "0010100100010100", 
        "0010100111101110", 
        "0010101011000100", 
        "0010101110010111", 
        "0010110001100111", 
        "0010110100110011", 
        "0010110111111011", 
        "0010111011000000", 
        "0010111110000010", 
        "0011000000111111", 
        "0011000011111001", 
        "0011000110101111", 
        "0011001001100010", 
        "0011001100010000", 
        "0011001110111010", 
        "0011010001100000", 
        "0011010100000011", 
        "0011010110100001", 
        "0011011000111011", 
        "0011011011010000", 
        "0011011101100010", 
        "0011011111101111", 
        "0011100001110111", 
        "0011100011111100", 
        "0011100101111100", 
        "0011100111110111", 
        "0011101001101110", 
        "0011101011100000", 
        "0011101101001110", 
        "0011101110110111", 
        "0011110000011011", 
        "0011110001111011", 
        "0011110011010110", 
        "0011110100101101", 
        "0011110101111110", 
        "0011110111001011", 
        "0011111000010011", 
        "0011111001010110", 
        "0011111010010100", 
        "0011111011001110", 
        "0011111100000010", 
        "0011111100110010", 
        "0011111101011101", 
        "0011111110000010", 
        "0011111110100011", 
        "0011111110111111", 
        "0011111111010110", 
        "0011111111101000", 
        "0011111111110101", 
        "0011111111111101", 
        "0011111111111111", 
        "0011111111111101", 
        "0011111111110110", 
        "0011111111101010", 
        "0011111111011001", 
        "0011111111000011", 
        "0011111110101001", 
        "0011111110001001", 
        "0011111101100100", 
        "0011111100111010", 
        "0011111100001011", 
        "0011111011011000", 
        "0011111010011111", 
        "0011111001100010", 
        "0011111000100000", 
        "0011110111011001", 
        "0011110110001101", 
        "0011110100111100", 
        "0011110011100110", 
        "0011110010001100", 
        "0011110000101101", 
        "0011101111001010", 
        "0011101101100001", 
        "0011101011110101", 
        "0011101010000011", 
        "0011101000001101", 
        "0011100110010010", 
        "0011100100010011", 
        "0011100010010000", 
        "0011100000001000", 
        "0011011101111100", 
        "0011011011101011", 
        "0011011001010110", 
        "0011010110111101", 
        "0011010100100000", 
        "0011010001111110", 
        "0011001111011001", 
        "0011001100101111", 
        "0011001010000010", 
        "0011000111010000", 
        "0011000100011011", 
        "0011000001100010", 
        "0010111110100101", 
        "0010111011100100", 
        "0010111000100000", 
        "0010110101011000", 
        "0010110010001100", 
        "0010101110111101", 
        "0010101011101011", 
        "0010101000010101", 
        "0010100100111100", 
        "0010100001100000", 
        "0010011110000001", 
        "0010011010011111", 
        "0010010110111001", 
        "0010010011010001", 
        "0010001111100110", 
        "0010001011111000", 
        "0010001000000111", 
        "0010000100010100", 
        "0010000000011110", 
        "0001111100100101", 
        "0001111000101010", 
        "0001110100101101", 
        "0001110000101110", 
        "0001101100101100", 
        "0001101000101000", 
        "0001100100100010", 
        "0001100000011010", 
        "0001011100010001", 
        "0001011000000101", 
        "0001010011111000", 
        "0001001111101001", 
        "0001001011011001", 
        "0001000111000111", 
        "0001000010110100", 
        "0000111110011111", 
        "0000111010001001", 
        "0000110101110011", 
        "0000110001011011", 
        "0000101101000010", 
        "0000101000101000", 
        "0000100100001101", 
        "0000011111110010", 
        "0000011011010110", 
        "0000010110111010", 
        "0000010010011101", 
        "0000001110000000", 
        "0000001001100010", 
        "0000000101000100", 
        "0000000000100111", 
        "0000000011110110", 
        "0000001000010100", 
        "0000001100110001", 
        "0000010001001111", 
        "0000010101101100", 
        "0000011010001000", 
        "0000011110100100", 
        "0000100011000000", 
        "0000100111011011", 
        "0000101011110101", 
        "0000110000001110", 
        "0000110100100110", 
        "0000111000111101", 
        "0000111101010011", 
        "0001000001101000", 
        "0001000101111100", 
        "0001001010001110", 
        "0001001110011111", 
        "0001010010101110", 
        "0001010110111100", 
        "0001011011001000", 
        "0001011111010010", 
        "0001100011011010", 
        "0001100111100001", 
        "0001101011100101", 
        "0001101111100111", 
        "0001110011100111", 
        "0001110111100101", 
        "0001111011100001", 
        "0001111111011010", 
        "0010000011010000", 
        "0010000111000101", 
        "0010001010110110", 
        "0010001110100101", 
        "0010010010010001", 
        "0010010101111010", 
        "0010011001100000", 
        "0010011101000011", 
        "0010100000100011", 
        "0010100100000000", 
        "0010100111011010", 
        "0010101010110001", 
        "0010101110000100", 
        "0010110001010100", 
        "0010110100100000", 
        "0010110111101001", 
        "0010111010101111", 
        "0010111101110000", 
        "0011000000101110", 
        "0011000011101001", 
        "0011000110011111", 
        "0011001001010001", 
        "0011001100000000", 
        "0011001110101011", 
        "0011010001010001", 
        "0011010011110100", 
        "0011010110010010", 
        "0011011000101101", 
        "0011011011000011", 
        "0011011101010100", 
        "0011011111100010", 
        "0011100001101011", 
        "0011100011110000", 
        "0011100101110000", 
        "0011100111101100", 
        "0011101001100011", 
        "0011101011010110", 
        "0011101101000100", 
        "0011101110101110", 
        "0011110000010010", 
        "0011110001110011", 
        "0011110011001110", 
        "0011110100100101", 
        "0011110101110111", 
        "0011110111000100", 
        "0011111000001101", 
        "0011111001010000", 
        "0011111010001111", 
        "0011111011001001", 
        "0011111011111110", 
        "0011111100101110", 
        "0011111101011001", 
        "0011111101111111", 
        "0011111110100000", 
        "0011111110111101", 
        "0011111111010100", 
        "0011111111100110", 
        "0011111111110100", 
        "0011111111111100"

    );

begin
    process(clk, angle)

    begin
        
        if clk'event and clk = '1' then
            if en = '1' then
                cos <= ROM(to_integer(unsigned(angle)));
            end if;
        end if;
    end process;


end syn;
