----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/06/2023 04:13:28 PM
-- Design Name: 
-- Module Name: RAM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with unsigned or unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity roms_tsp is
    Generic(
        WIDTH_D: positive;
        WIDTH_A: positive;
        DEPTH: positive
    );
    Port (
        clk: in std_logic;

        addr_i: in std_logic_vector(WIDTH_A-1 downto 0);
        data_o: out std_logic_vector(WIDTH_D-1 downto 0);

        en: in std_logic
    );
end roms_tsp;

architecture syn of roms_tsp is

    type rom_type is array(0 to DEPTH-1) of std_logic_vector(WIDTH_D-1 downto 0);
    signal ROM: rom_type :=(
        "0000001011001010",
        "0000100001011010",
        "0000110111011010",
        "0001001100111110",
        "0001100001111101",
        "0001110110001101",
        "0010001001100011",
        "0010011011110101",
        "0010101100111100",
        "0010111100101111",
        "0011001011000110",
        "0011010111111010",
        "0011100011000100",
        "0011101100100000",
        "0011110100001001",
        "0011111001111011",
        "0011111101110011",
        "0011111111110000",
        "0011111111110000",
        "0011111101110011",
        "0011111001111011",
        "0011110100001001",
        "0011101100100000",
        "0011100011000100",
        "0011010111111010",
        "0011001011000110",
        "0010111100101111",
        "0010101100111100",
        "0010011011110101",
        "0010001001100011",
        "0001110110001101",
        "0001100001111101",
        "0001001100111110",
        "0000110111011010",
        "0000100001011010",
        "0000001011001010",
        "0000001011001010",
        "0000100001011010",
        "0000110111011010",
        "0001001100111110",
        "0001100001111101",
        "0001110110001101",
        "0010001001100011",
        "0010011011110101",
        "0010101100111100",
        "0010111100101111",
        "0011001011000110",
        "0011010111111010",
        "0011100011000100",
        "0011101100100000",
        "0011110100001001",
        "0011111001111011",
        "0011111101110011",
        "0011111111110000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0011111101110011",
        "0011101100100000",
        "0011001011000110",
        "0010011011110101",
        "0001100001111101",
        "0000100001011010",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000100001011010",
        "0001100001111101",
        "0010011011110101",
        "0011001011000110",
        "0011101100100000",
        "0011111101110011",
        "0011111101110011",
        "0011101100100000",
        "0011001011000110",
        "0010011011110101",
        "0001100001111101",
        "0000100001011010",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000100001011010",
        "0001100001111101",
        "0010011011110101",
        "0011001011000110",
        "0011101100100000",
        "0011111101110011",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0100000000000000",
        "0011111111110000",
        "0011111101110011",
        "0011111001111011",
        "0011110100001001",
        "0011101100100000",
        "0011100011000100",
        "0011010111111010",
        "0011001011000110",
        "0010111100101111",
        "0010101100111100",
        "0010011011110101",
        "0010001001100011",
        "0001110110001101",
        "0001100001111101",
        "0001001100111110",
        "0000110111011010",
        "0000100001011010",
        "0000001011001010"
    );
begin
    process(clk, addr_i)
    begin
        if clk'event and clk = '1' then
            if en = '1' then
                data_o <= ROM(to_integer(unsigned(addr_i)));
            end if;
        end if;
    end process;

end syn;





















